library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

use work.common_types.all;

entity rr_arbiter_321 is
    generic (
        DWIDTH : natural := 39 -- data word width from requester FIFOs
    );
    port (
        -- Input from requesters 
        empty_in : std_logic_vector(0 to 31);    -- Empty signals from requester FIFOs
        valid_in : std_logic_vector(0 to 31);    -- Read valid signals from requester FIFOs
        data_in  : SlvArray(0 to 31)(DWIDTH-1 downto 0);         -- Read data from requester FIFOs
        -- Control inputs
        clk      : in std_logic;    -- 4x system clock (212.4 MHz)
        rst      : in std_logic;    -- synchronous, active high reset
        -- Outputs
        enable_out : out std_logic_vector(0 to 31);  -- Read enable signals sent to requester FIFOs
        data_out   : out std_logic_vector(DWIDTH-1 downto 0);   -- Data from granted requester, sent to event ring buffer
        valid_out  : out std_logic     -- sent to wr_enable of the event ring buffer alongside data_out
    );
end rr_arbiter_321;

architecture Behavioral of rr_arbiter_321 is

    type state is (s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_tx);
    signal present_state, next_state, buffer_state: state;
    -- Register the request and grant 
    signal request_reg, grant_reg : std_logic_vector(0 to 31);
    -- Store an integer to determine which of the inputs has been granted
    signal which_fifo : integer range 0 to 31;
    
begin

    -- Invert the empty signals from the FIFOs to act as the request register
    process(all)
    begin
        if rising_edge(clk) then
            request_reg <= not empty_in;
        end if;
    end process;
    
    -- Monitor the request register and issue grants based on round-robin arbitration.
    -- When a request is observed (a non-empty requester FIFO), a grant is issued and the 
    -- state moves to transmit, where a FIFO read is granted and the system waits for the 
    -- read valid flag from the FIFO. After the read valid flag is pulsed, the state machine
    -- moves to the buffered state and the process continues until there are no more requests.
    arbitrate : process(all)
    begin
        if rising_edge(clk) then
            if rst = '1' then 
                valid_out     <= '0';
                data_out      <= (others => '0');
                enable_out    <= (others => '0');
                buffer_state  <= s_0;
                next_state    <= s_0;
                present_state <= s_0;
                which_fifo    <= 0;
            else
                present_state <= next_state;
                case present_state is
                    when s_0 =>
                        valid_out <= '0';
                        if request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_1 =>
                        valid_out <= '0';
                        if request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_2 =>
                        valid_out <= '0';
                        if request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_3 =>
                        valid_out <= '0';
                        if request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_4 =>
                        valid_out <= '0';
                        if request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_5 =>
                        valid_out <= '0';
                        if request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_6 =>
                        valid_out <= '0';
                        if request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_7 =>
                        valid_out <= '0';
                        if request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_8 =>
                        valid_out <= '0';
                        if request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_9 =>
                        valid_out <= '0';
                        if request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_10 =>
                        valid_out <= '0';
                        if request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_11 =>
                        valid_out <= '0';
                        if request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_12 =>
                        valid_out <= '0';
                        if request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_13 =>
                        valid_out <= '0';
                        if request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_14 =>
                        valid_out <= '0';
                        if request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_15 =>
                        valid_out <= '0';
                        if request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_16 =>
                        valid_out <= '0';
                        if request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_17 =>
                        valid_out <= '0';
                        if request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_18 =>
                        valid_out <= '0';
                        if request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_19 =>
                        valid_out <= '0';
                        if request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_20 =>
                        valid_out <= '0';
                        if request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_21 =>
                        valid_out <= '0';
                        if request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_22 =>
                        valid_out <= '0';
                        if request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_23 =>
                        valid_out <= '0';
                        if request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_24 =>
                        valid_out <= '0';
                        if request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_25 =>
                        valid_out <= '0';
                        if request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_26 =>
                        valid_out <= '0';
                        if request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_27 =>
                        valid_out <= '0';
                        if request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_28 =>
                        valid_out <= '0';
                        if request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_29 =>
                        valid_out <= '0';
                        if request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_30 =>
                        valid_out <= '0';
                        if request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        elsif request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_31 =>
                        valid_out <= '0';
                        if request_reg(31) = '1' then
                            grant_reg    <= "00000000000000000000000000000001";
                            enable_out   <= "00000000000000000000000000000001";
                            which_fifo   <= 31;
                            next_state   <= s_tx;
                            buffer_state <= s_0;
                        elsif request_reg(0) = '1' then
                            grant_reg    <= "10000000000000000000000000000000";
                            enable_out   <= "10000000000000000000000000000000";
                            which_fifo   <= 0;
                            next_state   <= s_tx;
                            buffer_state <= s_1;
                        elsif request_reg(1) = '1' then
                            grant_reg    <= "01000000000000000000000000000000";
                            enable_out   <= "01000000000000000000000000000000";
                            which_fifo   <= 1;
                            next_state   <= s_tx;
                            buffer_state <= s_2;
                        elsif request_reg(2) = '1' then
                            grant_reg    <= "00100000000000000000000000000000";
                            enable_out   <= "00100000000000000000000000000000";
                            which_fifo   <= 2;
                            next_state   <= s_tx;
                            buffer_state <= s_3;
                        elsif request_reg(3) = '1' then
                            grant_reg    <= "00010000000000000000000000000000";
                            enable_out   <= "00010000000000000000000000000000";
                            which_fifo   <= 3;
                            next_state   <= s_tx;
                            buffer_state <= s_4;
                        elsif request_reg(4) = '1' then
                            grant_reg    <= "00001000000000000000000000000000";
                            enable_out   <= "00001000000000000000000000000000";
                            which_fifo   <= 4;
                            next_state   <= s_tx;
                            buffer_state <= s_5;
                        elsif request_reg(5) = '1' then
                            grant_reg    <= "00000100000000000000000000000000";
                            enable_out   <= "00000100000000000000000000000000";
                            which_fifo   <= 5;
                            next_state   <= s_tx;
                            buffer_state <= s_6;
                        elsif request_reg(6) = '1' then
                            grant_reg    <= "00000010000000000000000000000000";
                            enable_out   <= "00000010000000000000000000000000";
                            which_fifo   <= 6;
                            next_state   <= s_tx;
                            buffer_state <= s_7;
                        elsif request_reg(7) = '1' then
                            grant_reg    <= "00000001000000000000000000000000";
                            enable_out   <= "00000001000000000000000000000000";
                            which_fifo   <= 7;
                            next_state   <= s_tx;
                            buffer_state <= s_8;
                        elsif request_reg(8) = '1' then
                            grant_reg    <= "00000000100000000000000000000000";
                            enable_out   <= "00000000100000000000000000000000";
                            which_fifo   <= 8;
                            next_state   <= s_tx;
                            buffer_state <= s_9;
                        elsif request_reg(9) = '1' then
                            grant_reg    <= "00000000010000000000000000000000";
                            enable_out   <= "00000000010000000000000000000000";
                            which_fifo   <= 9;
                            next_state   <= s_tx;
                            buffer_state <= s_10;
                        elsif request_reg(10) = '1' then
                            grant_reg    <= "00000000001000000000000000000000";
                            enable_out   <= "00000000001000000000000000000000";
                            which_fifo   <= 10;
                            next_state   <= s_tx;
                            buffer_state <= s_11;
                        elsif request_reg(11) = '1' then
                            grant_reg    <= "00000000000100000000000000000000";
                            enable_out   <= "00000000000100000000000000000000";
                            which_fifo   <= 11;
                            next_state   <= s_tx;
                            buffer_state <= s_12;
                        elsif request_reg(12) = '1' then
                            grant_reg    <= "00000000000010000000000000000000";
                            enable_out   <= "00000000000010000000000000000000";
                            which_fifo   <= 12;
                            next_state   <= s_tx;
                            buffer_state <= s_13;
                        elsif request_reg(13) = '1' then
                            grant_reg    <= "00000000000001000000000000000000";
                            enable_out   <= "00000000000001000000000000000000";
                            which_fifo   <= 13;
                            next_state   <= s_tx;
                            buffer_state <= s_14;
                        elsif request_reg(14) = '1' then
                            grant_reg    <= "00000000000000100000000000000000";
                            enable_out   <= "00000000000000100000000000000000";
                            which_fifo   <= 14;
                            next_state   <= s_tx;
                            buffer_state <= s_15;
                        elsif request_reg(15) = '1' then
                            grant_reg    <= "00000000000000010000000000000000";
                            enable_out   <= "00000000000000010000000000000000";
                            which_fifo   <= 15;
                            next_state   <= s_tx;
                            buffer_state <= s_16;
                        elsif request_reg(16) = '1' then
                            grant_reg    <= "00000000000000001000000000000000";
                            enable_out   <= "00000000000000001000000000000000";
                            which_fifo   <= 16;
                            next_state   <= s_tx;
                            buffer_state <= s_17;
                        elsif request_reg(17) = '1' then
                            grant_reg    <= "00000000000000000100000000000000";
                            enable_out   <= "00000000000000000100000000000000";
                            which_fifo   <= 17;
                            next_state   <= s_tx;
                            buffer_state <= s_18;
                        elsif request_reg(18) = '1' then
                            grant_reg    <= "00000000000000000010000000000000";
                            enable_out   <= "00000000000000000010000000000000";
                            which_fifo   <= 18;
                            next_state   <= s_tx;
                            buffer_state <= s_19;
                        elsif request_reg(19) = '1' then
                            grant_reg    <= "00000000000000000001000000000000";
                            enable_out   <= "00000000000000000001000000000000";
                            which_fifo   <= 19;
                            next_state   <= s_tx;
                            buffer_state <= s_20;
                        elsif request_reg(20) = '1' then
                            grant_reg    <= "00000000000000000000100000000000";
                            enable_out   <= "00000000000000000000100000000000";
                            which_fifo   <= 20;
                            next_state   <= s_tx;
                            buffer_state <= s_21;
                        elsif request_reg(21) = '1' then
                            grant_reg    <= "00000000000000000000010000000000";
                            enable_out   <= "00000000000000000000010000000000";
                            which_fifo   <= 21;
                            next_state   <= s_tx;
                            buffer_state <= s_22;
                        elsif request_reg(22) = '1' then
                            grant_reg    <= "00000000000000000000001000000000";
                            enable_out   <= "00000000000000000000001000000000";
                            which_fifo   <= 22;
                            next_state   <= s_tx;
                            buffer_state <= s_23;
                        elsif request_reg(23) = '1' then
                            grant_reg    <= "00000000000000000000000100000000";
                            enable_out   <= "00000000000000000000000100000000";
                            which_fifo   <= 23;
                            next_state   <= s_tx;
                            buffer_state <= s_24;
                        elsif request_reg(24) = '1' then
                            grant_reg    <= "00000000000000000000000010000000";
                            enable_out   <= "00000000000000000000000010000000";
                            which_fifo   <= 24;
                            next_state   <= s_tx;
                            buffer_state <= s_25;
                        elsif request_reg(25) = '1' then
                            grant_reg    <= "00000000000000000000000001000000";
                            enable_out   <= "00000000000000000000000001000000";
                            which_fifo   <= 25;
                            next_state   <= s_tx;
                            buffer_state <= s_26;
                        elsif request_reg(26) = '1' then
                            grant_reg    <= "00000000000000000000000000100000";
                            enable_out   <= "00000000000000000000000000100000";
                            which_fifo   <= 26;
                            next_state   <= s_tx;
                            buffer_state <= s_27;
                        elsif request_reg(27) = '1' then
                            grant_reg    <= "00000000000000000000000000010000";
                            enable_out   <= "00000000000000000000000000010000";
                            which_fifo   <= 27;
                            next_state   <= s_tx;
                            buffer_state <= s_28;
                        elsif request_reg(28) = '1' then
                            grant_reg    <= "00000000000000000000000000001000";
                            enable_out   <= "00000000000000000000000000001000";
                            which_fifo   <= 28;
                            next_state   <= s_tx;
                            buffer_state <= s_29;
                        elsif request_reg(29) = '1' then
                            grant_reg    <= "00000000000000000000000000000100";
                            enable_out   <= "00000000000000000000000000000100";
                            which_fifo   <= 29;
                            next_state   <= s_tx;
                            buffer_state <= s_30;
                        elsif request_reg(30) = '1' then
                            grant_reg    <= "00000000000000000000000000000010";
                            enable_out   <= "00000000000000000000000000000010";
                            which_fifo   <= 30;
                            next_state   <= s_tx;
                            buffer_state <= s_31;
                        else
                            grant_reg    <= (others => '0');
                            enable_out   <= (others => '0');
                            which_fifo   <= 0;
                            next_state   <= s_0;
                            buffer_state <= s_0;
                        end if;
                    when s_tx =>
                        -- disable the read_enable so it's only high for one clock period (avoids losing data in the FIFO if there are multiple hits)
                        enable_out(which_fifo) <= '0';
                        -- Tie the data output to the read data of the granted FIFO requester
                        data_out <= data_in(which_fifo);
                        valid_out <= '1';
                        -- wait for the FIFO to return the valid read flag before moving to next (buffered) state
                        if valid_in(which_fifo) = '1' then 
                            -- The FIFO has successfully read out
                            next_state <= buffer_state; -- move to next state in round robin
                        end if;
                    when others => 
                        grant_reg    <= (others => '0');
                        enable_out   <= (others => '0');
                        which_fifo   <= 0;
                        next_state   <= s_0;
                        buffer_state <= s_0;
                end case;
            end if;
        end if;
    end process arbitrate;

end Behavioral;
